//Provided HDMI_Text_controller_v1_0 for HDMI AXI4 IP 
//Fall 2024 Distribution

//Modified 3/10/24 by Zuofu
//Updated 11/18/24 by Zuofu


`timescale 1 ns / 1 ps

module little_alchemy_controller_v1_0 #
(
    // Parameters of Axi Slave Bus Interface S00_AXI
    // Modify parameters as necessary for access of full VRAM range

    parameter integer C_AXI_DATA_WIDTH	= 32,
    parameter integer C_AXI_ADDR_WIDTH	= 16 
)
(
    input logic [31:0] mouse_gpio,
    // Users to add ports here

    output logic hdmi_clk_n,
    output logic hdmi_clk_p,
    output logic [2:0] hdmi_tx_n,
    output logic [2:0] hdmi_tx_p,

    // User ports ends
    // Do not modify the ports beyond this line


    // Ports of Axi Slave Bus Interface AXI
    input logic  axi_aclk,
    input logic  axi_aresetn,
    input logic [C_AXI_ADDR_WIDTH-1 : 0] axi_awaddr,
    input logic [2 : 0] axi_awprot,
    input logic  axi_awvalid,
    output logic  axi_awready,
    input logic [C_AXI_DATA_WIDTH-1 : 0] axi_wdata,
    input logic [(C_AXI_DATA_WIDTH/8)-1 : 0] axi_wstrb,
    input logic  axi_wvalid,
    output logic  axi_wready,
    output logic [1 : 0] axi_bresp,
    output logic  axi_bvalid,
    input logic  axi_bready,
    input logic [C_AXI_ADDR_WIDTH-1 : 0] axi_araddr,
    input logic [2 : 0] axi_arprot,
    input logic  axi_arvalid,
    output logic  axi_arready,
    output logic [C_AXI_DATA_WIDTH-1 : 0] axi_rdata,
    output logic [1 : 0] axi_rresp,
    output logic  axi_rvalid,
    input logic  axi_rready
);

//additional logic variables as necessary to support VGA, and HDMI modules.
    logic clk_25MHz, clk_125MHz;
    logic locked;
    logic [9:0] drawX, drawY;
    
    logic hsync, vsync, vde;
    logic [7:0] red, green, blue;
    logic [17:0] pixel_addr;
    logic [13:0] char_addr;
    logic [7:0]  char_idx;
    
    logic [7:0] pixel_color_idx;
    
    
    logic reset_ah;
    
    logic [C_AXI_DATA_WIDTH - 1:0] frame_cnt;
    assign reset_ah = ~axi_aresetn;
    logic [9:0] Mouse_X, Mouse_Y;
    logic signed [7:0] Mouse_XDiff, Mouse_YDiff;
    logic [7:0] Scroll_Diff;
    logic [7:0] Buttons;
    logic [9:0] MouseElementIdx;
    
    logic [9:0]  bram_addra, bram_addrb;
    logic [31:0]  bram_dina, bram_dinb;
    logic [0:0]   bram_wea;
    logic [31:0]  bram_douta, bram_doutb;
    
    logic [4:0]   MenuSlotIdx;
    logic [9:0]   MenuElementIdx;
    logic         ScreenMode;
    logic [9:0]   NewElement;
    
    
    
    assign Buttons = mouse_gpio[7:0];
    assign Mouse_XDiff = mouse_gpio[15:8];
    assign Mouse_YDiff = mouse_gpio[23:16];
    assign Scroll_Diff = mouse_gpio[31:24];
    
// Instantiation of Axi Bus Interface AXI
little_alchemy_controller_v1_0_AXI # ( 
    .C_S_AXI_DATA_WIDTH(C_AXI_DATA_WIDTH),
    .C_S_AXI_ADDR_WIDTH(C_AXI_ADDR_WIDTH)
) little_alchemy_controller_v1_0_AXI_inst (
    .frame_cnt(frame_cnt),
    .cur_draw_x(drawX),
    .cur_draw_y(drawY),
    .Mouse_X(Mouse_X),
    .Mouse_Y(Mouse_Y),
    .MenuSlotIdx(MenuSlotIdx),
    .MenuElementIdx(MenuElementIdx),
    .bram_douta(bram_douta),
    .bram_addra(bram_addra),
    .bram_dina(bram_dina),
    .bram_wea(bram_wea),
    .Mouse_Element(MouseElementIdx),
    .NewElement(NewElement),
    .ScreenMode(ScreenMode),
    .S_AXI_ACLK(axi_aclk),
    .S_AXI_ARESETN(axi_aresetn),
    .S_AXI_AWADDR(axi_awaddr),
    .S_AXI_AWPROT(axi_awprot),
    .S_AXI_AWVALID(axi_awvalid),
    .S_AXI_AWREADY(axi_awready),
    .S_AXI_WDATA(axi_wdata),
    .S_AXI_WSTRB(axi_wstrb),
    .S_AXI_WVALID(axi_wvalid),
    .S_AXI_WREADY(axi_wready),
    .S_AXI_BRESP(axi_bresp),
    .S_AXI_BVALID(axi_bvalid),
    .S_AXI_BREADY(axi_bready),
    .S_AXI_ARADDR(axi_araddr),
    .S_AXI_ARPROT(axi_arprot),
    .S_AXI_ARVALID(axi_arvalid),
    .S_AXI_ARREADY(axi_arready),
    .S_AXI_RDATA(axi_rdata),
    .S_AXI_RRESP(axi_rresp),
    .S_AXI_RVALID(axi_rvalid),
    .S_AXI_RREADY(axi_rready)
);


//Instiante clocking wizard, VGA sync generator modules, and VGA-HDMI IP here. For a hint, refer to the provided
//top-level from the previous lab. You should get the IP to generate a valid HDMI signal (e.g. blue screen or gradient)
//prior to working on the text drawing.

// User logic ends
    //clock wizard configured with a 1x and 5x clock for HDMI
    clk_wiz_0 clk_wiz (
        .clk_out1(clk_25MHz),
        .clk_out2(clk_125MHz),
        .reset(reset_ah),
        .locked(locked),
        .clk_in1(axi_aclk)
    );
    
    //VGA Sync signal generator
    vga_controller vga (
        .pixel_clk(clk_25MHz),
        .reset(reset_ah),
        .hs(hsync),
        .vs(vsync),
        .active_nblank(vde),
        .drawX(drawX),
        .drawY(drawY)
    );    

    //Real Digital VGA to HDMI converter
    hdmi_tx_0 vga_to_hdmi (
        //Clocking and Reset
        .pix_clk(clk_25MHz),
        .pix_clkx5(clk_125MHz),
        .pix_clk_locked(locked),
        .rst(reset_ah),
        //Color and Sync Signals
        .red(red),
        .green(green),
        .blue(blue),
        .hsync(hsync),
        .vsync(vsync),
        .vde(vde),
        
        //aux Data (unused)
        .aux0_din(4'b0),
        .aux1_din(4'b0),
        .aux2_din(4'b0),
        .ade(1'b0),
        
        //Differential outputs
        .TMDS_CLK_P(hdmi_clk_p),          
        .TMDS_CLK_N(hdmi_clk_n),          
        .TMDS_DATA_P(hdmi_tx_p),         
        .TMDS_DATA_N(hdmi_tx_n)          
    );

    
    //Color Mapper Module   
    color_mapper color_instance(
        .ScreenMode(ScreenMode),
        .DrawX(drawX),
        .DrawY(drawY),
        .MouseX(Mouse_X),
        .MouseY(Mouse_Y),
        .CharAddress(char_addr),
        .CharIdx(char_idx),
        .MouseElementIdx(MouseElementIdx),
        .WorkspaceElementIdx(bram_doutb),
        .MenuElementIdx(MenuElementIdx),
        .NewElement(NewElement),
        .PixelAddress(pixel_addr),
        .PaletteIdx(pixel_color_idx),
        .WorkspaceSlotIdx(bram_addrb),
        .MenuSlotIdx(MenuSlotIdx),
        .Red(red),
        .Green(green),
        .Blue(blue)
    );
    
    frame_counter frame_counter_inst(
    .Reset(reset_ah),
    .frame_clk(~vsync), 
    .frame_cnt(frame_cnt)
    );
    
    mouse mouse_inst (
    .Reset(reset_ah),
    .frame_clk(~vsync),
    .Mouse_XDiff(Mouse_XDiff),
    .Mouse_YDiff(Mouse_YDiff),
    .Buttons(Buttons),
    .Mouse_X(Mouse_X),
    .Mouse_Y(Mouse_Y)
    );
    
    little_alchemy_graphics_rom graphics_rom(
        .clka(axi_aclk),
        .addra(pixel_addr),
        .douta(pixel_color_idx)
    ); 
    element_text_rom little_alchemy_text_rom(
        .clka(axi_aclk),
        .addra(char_addr),
        .douta(char_idx)
    ); 
    
    workspace_blk_mem workspace_bram (
        .addra	(bram_addra),
        .clka	(axi_aclk),
        .dina	(bram_dina),
        .wea	(bram_wea),
        .douta	(bram_douta),
        .addrb	(bram_addrb),
        .clkb	(axi_aclk),
        .dinb	(0),
        .web	(0),
        .doutb	(bram_doutb)
    );
    

endmodule
